V1 1 0 1
R1 1 0 1

.control
    .op
.end
