V1 1 0 1
R1 1 2 1
R2 2 0 1

.control
    .op
.end
